module ctr (
	input	wire	clk,
	input 	wire	rst
);

endmodule